library ieee;
use ieee.std_logic_1164.all;

entity aes_sbox is
    port (
        datai : in  std_logic_vector(7 downto 0);
        datao : out std_logic_vector(7 downto 0)
    );
end entity;

architecture rtl of aes_sbox is
    signal u0   : std_logic;
    signal u1   : std_logic;
    signal u2   : std_logic;
    signal u3   : std_logic;
    signal u4   : std_logic;
    signal u5   : std_logic;
    signal u6   : std_logic;
    signal u7   : std_logic;

    signal y14  : std_logic;
    signal y13  : std_logic;
    signal y9   : std_logic;
    signal y8   : std_logic;
    signal t0   : std_logic;
    signal y1   : std_logic;
    signal y4   : std_logic;
    signal y12  : std_logic;
    signal y2   : std_logic;
    signal y5   : std_logic;
    signal y3   : std_logic;
    signal t1   : std_logic;
    signal y15  : std_logic;
    signal y20  : std_logic;
    signal y6   : std_logic;
    signal y10  : std_logic;
    signal y11  : std_logic;
    signal y7   : std_logic;
    signal y17  : std_logic;
    signal y19  : std_logic;
    signal y16  : std_logic;
    signal y21  : std_logic;
    signal y18  : std_logic;
    signal t2   : std_logic;
    signal t3   : std_logic;
    signal t4   : std_logic;
    signal t5   : std_logic;
    signal t6   : std_logic;
    signal t7   : std_logic;
    signal t8   : std_logic;
    signal t9   : std_logic;
    signal t10  : std_logic;
    signal t11  : std_logic;
    signal t12  : std_logic;
    signal t13  : std_logic;
    signal t14  : std_logic;
    signal t15  : std_logic;
    signal t16  : std_logic;
    signal t17  : std_logic;
    signal t18  : std_logic;
    signal t19  : std_logic;
    signal t20  : std_logic;
    signal t21  : std_logic;
    signal t22  : std_logic;
    signal t23  : std_logic;
    signal t24  : std_logic;
    signal t25  : std_logic;
    signal t26  : std_logic;
    signal t27  : std_logic;
    signal t28  : std_logic;
    signal t29  : std_logic;
    signal t30  : std_logic;
    signal t31  : std_logic;
    signal t32  : std_logic;
    signal t33  : std_logic;
    signal t34  : std_logic;
    signal t35  : std_logic;
    signal t36  : std_logic;
    signal t37  : std_logic;
    signal t38  : std_logic;
    signal t39  : std_logic;
    signal t40  : std_logic;
    signal t41  : std_logic;
    signal t42  : std_logic;
    signal t43  : std_logic;
    signal t44  : std_logic;
    signal t45  : std_logic;
    signal z0   : std_logic;
    signal z1   : std_logic;
    signal z2   : std_logic;
    signal z3   : std_logic;
    signal z4   : std_logic;
    signal z5   : std_logic;
    signal z6   : std_logic;
    signal z7   : std_logic;
    signal z8   : std_logic;
    signal z9   : std_logic;
    signal z10  : std_logic;
    signal z11  : std_logic;
    signal z12  : std_logic;
    signal z13  : std_logic;
    signal z14  : std_logic;
    signal z15  : std_logic;
    signal z16  : std_logic;
    signal z17  : std_logic;
    signal tc1  : std_logic;
    signal tc2  : std_logic;
    signal tc3  : std_logic;
    signal tc4  : std_logic;
    signal tc5  : std_logic;
    signal tc6  : std_logic;
    signal tc7  : std_logic;
    signal tc8  : std_logic;
    signal tc9  : std_logic;
    signal tc10 : std_logic;
    signal tc11 : std_logic;
    signal tc12 : std_logic;
    signal tc13 : std_logic;
    signal tc14 : std_logic;
    signal tc16 : std_logic;
    signal tc17 : std_logic;
    signal tc18 : std_logic;
    signal tc20 : std_logic;
    signal tc21 : std_logic;
    signal tc26 : std_logic;

    signal s0   : std_logic;
    signal s1   : std_logic;
    signal s2   : std_logic;
    signal s3   : std_logic;
    signal s4   : std_logic;
    signal s5   : std_logic;
    signal s6   : std_logic;
    signal s7   : std_logic;
begin
    u0       <= datai(7);
    u1       <= datai(6);
    u2       <= datai(5);
    u3       <= datai(4);
    u4       <= datai(3);
    u5       <= datai(2);
    u6       <= datai(1);
    u7       <= datai(0);

    y14      <= u3   xor  u5;
    y13      <= u0   xor  u6;
    y9       <= u0   xor  u3;
    y8       <= u0   xor  u5;
    t0       <= u1   xor  u2;
    y1       <= t0   xor  u7;
    y4       <= y1   xor  u3;
    y12      <= y13  xor  y14;
    y2       <= y1   xor  u0;
    y5       <= y1   xor  u6;
    y3       <= y5   xor  y8;
    t1       <= u4   xor  y12;
    y15      <= t1   xor  u5;
    y20      <= t1   xor  u1;
    y6       <= y15  xor  u7;
    y10      <= y15  xor  t0;
    y11      <= y20  xor  y9;
    y7       <= u7   xor  y11;
    y17      <= y10  xor  y11;
    y19      <= y10  xor  y8;
    y16      <= t0   xor  y11;
    y21      <= y13  xor  y16;
    y18      <= u0   xor  y16;
    t2       <= y12  and  y15;
    t3       <= y3   and  y6;
    t4       <= t3   xor  t2;
    t5       <= y4   and  u7;
    t6       <= t5   xor  t2;
    t7       <= y13  and  y16;
    t8       <= y5   and  y1;
    t9       <= t8   xor  t7;
    t10      <= y2   and  y7;
    t11      <= t10  xor  t7;
    t12      <= y9   and  y11;
    t13      <= y14  and  y17;
    t14      <= t13  xor  t12;
    t15      <= y8   and  y10;
    t16      <= t15  xor  t12;
    t17      <= t4   xor  y20;
    t18      <= t6   xor  t16;
    t19      <= t9   xor  t14;
    t20      <= t11  xor  t16;
    t21      <= t17  xor  t14;
    t22      <= t18  xor  y19;
    t23      <= t19  xor  y21;
    t24      <= t20  xor  y18;
    t25      <= t21  xor  t22;
    t26      <= t21  and  t23;
    t27      <= t24  xor  t26;
    t28      <= t25  and  t27;
    t29      <= t28  xor  t22;
    t30      <= t23  xor  t24;
    t31      <= t22  xor  t26;
    t32      <= t31  and  t30;
    t33      <= t32  xor  t24;
    t34      <= t23  xor  t33;
    t35      <= t27  xor  t33;
    t36      <= t24  and  t35;
    t37      <= t36  xor  t34;
    t38      <= t27  xor  t36;
    t39      <= t29  and  t38;
    t40      <= t25  xor  t39;
    t41      <= t40  xor  t37;
    t42      <= t29  xor  t33;
    t43      <= t29  xor  t40;
    t44      <= t33  xor  t37;
    t45      <= t42  xor  t41;
    z0       <= t44  and  y15;
    z1       <= t37  and  y6;
    z2       <= t33  and  u7;
    z3       <= t43  and  y16;
    z4       <= t40  and  y1;
    z5       <= t29  and  y7;
    z6       <= t42  and  y11;
    z7       <= t45  and  y17;
    z8       <= t41  and  y10;
    z9       <= t44  and  y12;
    z10      <= t37  and  y3;
    z11      <= t33  and  y4;
    z12      <= t43  and  y13;
    z13      <= t40  and  y5;
    z14      <= t29  and  y2;
    z15      <= t42  and  y9;
    z16      <= t45  and  y14;
    z17      <= t41  and  y8;
    tc1      <= z15  xor  z16;
    tc2      <= z10  xor  tc1;
    tc3      <= z9   xor  tc2;
    tc4      <= z0   xor  z2;
    tc5      <= z1   xor  z0;
    tc6      <= z3   xor  z4;
    tc7      <= z12  xor  tc4;
    tc8      <= z7   xor  tc6;
    tc9      <= z8   xor  tc7;
    tc10     <= tc8  xor  tc9;
    tc11     <= tc6  xor  tc5;
    tc12     <= z3   xor  z5;
    tc13     <= z13  xor  tc1;
    tc14     <= tc4  xor  tc12;
    tc16     <= z6   xor  tc8;
    tc17     <= z14  xor  tc10;
    tc18     <= tc13 xor  tc14;
    tc20     <= z15  xor  tc16;
    tc21     <= tc2  xor  z11;
    tc26     <= tc17 xor  tc20;
    s3       <= tc3  xor  tc11;
    s7       <= z12  xnor tc18;
    s0       <= tc3  xor  tc16;
    s6       <= tc10 xnor tc18;
    s4       <= tc14 xor  s3;
    s1       <= s3   xnor tc16;
    s2       <= tc26 xnor z17;
    s5       <= tc21 xor  tc17;

    datao(7) <= s0;
    datao(6) <= s1;
    datao(5) <= s2;
    datao(4) <= s3;
    datao(3) <= s4;
    datao(2) <= s5;
    datao(1) <= s6;
    datao(0) <= s7;
end architecture rtl;
